module PU_tb;

endmodule
