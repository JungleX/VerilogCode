`define CTRL_WIDTH   16