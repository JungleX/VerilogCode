`define CTRL_WIDTH   30