`include "dw_params.vh"

module stratix_wrapper #(
	parameter DATA_WIDTH     = 16,
	parameter WEIGHT_WIDTH   = 16,
	parameter NUM_PE         = 8,
	parameter NUM_PU         = 150
)
(
	input wire         global_reset
);

wire locked;


endmodule
