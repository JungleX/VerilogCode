

module PU 
#(
	
	parameter integer OP_WIDTH        = 16,
	
	parameter integer NUM_PE          = 4




















)(
	input wire                               clk,
	input wire                               reset,
	
	input wire                               lrn_enable,
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	input wire [ DATA_IN_WIDTH  -1 : 0 ]    vecgen_wr_data
	
	
	
	
	
	
	
	
	
	
	
	
	
);




localparam integer DATA_IN_WIDTH     = OP_WIDTH * NUM_PE;









genvar i;




endmodule
