`timescale 1ns / 1ps

`include "CNN_Parameter.vh"

module CNNFSM(
    //input clk_p,
    //input clk_n,
    input rst,
    input clk,
    input transmission_start,
    
    output reg stop,
    output reg [7:0] led 
    );

	/*wire clk;

    IBUFDS #(
        .DIFF_TERM("FALSE"),
        .IBUF_LOW_PWR("TRUE"),
        .IOSTANDARD("DEFAULT")
         )IBUFDS_inst(
        .O(clk),
        .I(clk_p),
        .IB(clk_n)
    );*/

	reg lp_rst;

	reg [3:0] layer_type; // 0: prepare init feature map and weight data; 1:conv; 2:pool; 3:fc; 9: finish, done
	reg [3:0] pre_layer_type;

	reg [`LAYER_NUM_WIDTH - 1:0] layer_num;

	// data init and data update
	wire [`PARA_X*`POOL_SIZE*`PARA_Y*`DATA_WIDTH - 1:0] init_fm_data;
	wire [`WRITE_ADDR_WIDTH - 1:0] write_fm_data_addr;
	wire init_fm_data_done; // feature map data transmission, 0: not ready; 1: ready

	wire [`PARA_Y*`PARA_KERNEL*`DATA_WIDTH - 1:0] weight_data;
	wire [`WEIGHT_WRITE_ADDR_WIDTH*`PARA_KERNEL - 1:0] write_weight_data_addr;
	wire weight_data_done; // weight data transmission, 0: not ready; 1: ready

	// common configuration
	reg [`FM_SIZE_WIDTH - 1:0] fm_size;
	reg [`KERNEL_NUM_WIDTH - 1:0] fm_depth;
	reg [`FM_SIZE_WIDTH - 1:0] fm_total_size;

	reg [`FM_SIZE_WIDTH - 1:0] fm_size_out; // include padding
	reg [`PADDING_NUM_WIDTH - 1:0] padding_out;

	// conv
	reg [`KERNEL_NUM_WIDTH - 1:0] kernel_num; // fm_depth_out
	reg [`KERNEL_SIZE_WIDTH - 1:0] kernel_size;

	// pool
	reg pool_type; // 0: max pool; 1: avg pool
	reg [`POOL_SIZE_WIDTH - 1:0] pool_win_size; 

	// activation
	reg [1:0] activation; // 0: none; 1: ReLU. current just none or ReLU

	wire update_weight_ram; // 0: not update; 1: update
	wire [`WEIGHT_WRITE_ADDR_WIDTH - 1:0] update_weight_ram_addr;

	wire init_fm_ram_ready; // 0: not ready; 1: ready
	wire init_weight_ram_ready; // 0: not ready; 1: ready
	wire layer_ready;

	wire [`DATA_WIDTH - 1:0] test_data; // for debug
	// ======== Begin: layer ========
	LayerParaScaleFloat16 LP(
		.clk(clk),
		.rst(lp_rst),

		.layer_type(layer_type), // 0: prepare init feature map and weight data; 1:conv; 2:pool; 3:fc; 9: finish, done
		.pre_layer_type(pre_layer_type),

		.layer_num(layer_num),

		// data init and data update
		.init_fm_data(init_fm_data),
		.write_fm_data_addr(write_fm_data_addr),
		.init_fm_data_done(init_fm_data_done), // feature map data transmission, 0: not ready; 1: ready

		.weight_data(weight_data),
		.write_weight_data_addr(write_weight_data_addr),
		.weight_data_done(weight_data_done), // weight data transmission, 0: not ready; 1: ready

		// common configuration
		.fm_size(fm_size),
		.fm_depth(fm_depth),
		.fm_total_size(fm_total_size),

		.fm_size_out(fm_size_out), // include padding
		.padding_out(padding_out),

		// conv
		.kernel_num(kernel_num), // fm_depth_out
		.kernel_size(kernel_size),

		// pool
		.pool_type(pool_type), // 0: max pool; 1: avg pool
		.pool_win_size(pool_win_size), 

		// activation
		.activation(activation), // 0: none; 1: ReLU. current just none or ReLU

		.update_weight_ram(update_weight_ram), // 0: not update; 1: update
		.update_weight_ram_addr(update_weight_ram_addr),

		.init_fm_ram_ready(init_fm_ram_ready), // 0: not ready; 1: ready
		.init_weight_ram_ready(init_weight_ram_ready), // 0: not ready; 1: ready
		.layer_ready(layer_ready),

		.test_data(test_data)
    );
	// ======== End: layer ========

	reg dt_rst;

	reg [`WRITE_ADDR_WIDTH - 1:0] write_fm_num;

	reg [`KERNEL_NUM_WIDTH - 1:0] kernel_num_count;
    reg [`WEIGHT_READ_ADDR_WIDTH - 1:0] write_weight_num;
    reg [`WEIGHT_READ_ADDR_WIDTH - 1:0] next_write_weight_num;
	// ======== Begin: data ========
	DataTransFloat16 DT(
    	.clk(clk),
    	.rst(dt_rst),
    
    	.layer_type(layer_type),
    	.layer_num(layer_num),

    	.write_fm_num(write_fm_num),

    	.kernel_num_count(kernel_num_count),
    	.write_weight_num(write_weight_num),
    	.next_write_weight_num(next_write_weight_num),
    
    	.update_weight_ram(update_weight_ram), // 0: not update; 1: update
    	.update_weight_ram_addr(update_weight_ram_addr),
    
    	.init_fm_ram_ready(init_fm_ram_ready), // 0: not ready; 1: ready
    	.init_weight_ram_ready(init_weight_ram_ready), // 0: not ready; 1: ready
    
    	.init_fm_data(init_fm_data),
    	.write_fm_data_addr(write_fm_data_addr),
    	.init_fm_data_done(init_fm_data_done),
    
    	.weight_data(weight_data),
    	.write_weight_data_addr(write_weight_data_addr),
    	.weight_data_done(weight_data_done) // weight data transmission, 0: not ready; 1: ready
    );
	// ======== End: data ========

	reg workstate;
	reg [23:0] clk_cnt;
	reg [26:0] output_cnt;
	//reg [8:0] output_cnt;

	/*always @(transmission_start or rst or stop) 
    	workstate <= transmission_start & (rst) & (~stop);*/
    	
    always @(posedge clk or negedge rst) begin
    if (rst) workstate <= transmission_start;
    else if (!rst) workstate <= 0;
    end
    
    /*always @(posedge clk or negedge rst) begin
    if (!rst) stop <= 1'b0;
    else stop <= stop_cnt[30];
    end*/
    

    reg layer_delay;
	always @(posedge clk) 
    	layer_delay <= layer_ready;

    reg init_done;
    
    always @(posedge clk or negedge rst) begin
        if (!rst) stop <= 1'b0;
        else if (layer_type == 9) stop <= 1;
    end
                
    always @(posedge clk or negedge rst) begin
        if (!rst) clk_cnt <= 0;
        else if (workstate && !stop) clk_cnt <= clk_cnt + 1;
    end
        
    always @(posedge clk or negedge rst)
    if (!rst) output_cnt <= 0;
    else if(stop) output_cnt <= output_cnt + 1;
        
    always @(posedge clk)
        case (output_cnt[26:25])
        //case (output_cnt[8:7])
        2'b00:led <= 8'b0;
        2'b01:led <= clk_cnt[23:16];
        2'b10:led <= clk_cnt[15:8];
        2'b11:led <= clk_cnt[7:0];
        endcase

	always @(posedge clk or negedge rst) begin
		if (!rst) begin
			lp_rst <= 0;
			dt_rst <= 0;

			layer_type	<= 0;
			layer_num	<= 0;

			init_done			<= 0;
			write_fm_num		<= 0;
			write_weight_num	<= 0;
			next_write_weight_num <= 0;
			kernel_num_count	<= 0;
			
		end
		else begin
			if (workstate) begin
				if (init_done == 0) begin 
					layer_type		<= 0; 
			        layer_num		<= 0;

			        lp_rst			<= 1;
			        
			        dt_rst			<= 1;
			        
			        //write_fm_num	<= 12; // fm size: 8, depth: 2; [8/3] * [8/(2*3)] * 2 = 3 * 2 * 2 = 12
			        //write_weight_num<= 12; // kernel_size: 3; depth: 2; 3 * 3 * 2 * 2 / 3 = 12

			        // write_fm_num = [fm_size / `PARA_X] * [fm_size / (`POOL_SIZE * `PARA_Y)] * depth
			        // each ram save [fm_size / `PARA_X] line, each line write [fm_size / (`POOL_SIZE * `PARA_Y)] times
			        write_fm_num	<= ((28+`PARA_X-1)/`PARA_X) * ((28+(2*`PARA_Y)-1)/(2*`PARA_Y)) * 512; //25600; // fm size: 28, depth: 512; [28/3] * [28/(2*3)] * 512 = 10 * 5 * 512 = 25600
			        // write_weight_num = kernel_size * kernel_size * depth * 2 / `PARA_Y
			        write_weight_num<= (9216+`PARA_Y-1)/`PARA_Y; //3072; // kernel_size: 3; depth: 512; 3 * 3 * 512 * 2 / 3 = 3072; 3*3*512*2 = 9216
				end

				if ((layer_ready) && (~layer_delay)) begin // pre layer is ready, go to new layer
					init_done	<= 1;

					layer_num <= layer_num + 1;
			        case (layer_num + 1)
			            1: 
			            	begin 
			            		layer_type	<= 1; // conv
			        			activation	<= 1;

			        			fm_size		<= 28;
						        fm_depth	<= 4;  // 512 todo
						        fm_size_out <= 28; // including padding
						        padding_out <= 1;

						        kernel_num  <= 8; // 512 todo
						        kernel_size <= 3;

						        kernel_num_count <= 8 - `PARA_KERNEL*2; // 8 - `PARA_KERNEL*2 = 4 // 512 - `PARA_KERNEL*2 = 508 todo
						        write_weight_num <= (36+`PARA_Y-1)/`PARA_Y; // 3*3 * 4 = 36 // (4608+`PARA_Y-1)/`PARA_Y; 3*3 * 512 = 4608
						        next_write_weight_num <= (72+`PARA_Y-1)/`PARA_Y; //  3*3 * 8 = 72 // (4608+`PARA_Y-1)/`PARA_Y; 3*3 * 512 = 4608
			            	end
			            2:
			            	begin 
			            		layer_type		<= 2; // pool
			        			pool_type		<= 0;

						        pool_win_size	<= `POOL_SIZE;

						        fm_size 		<= 28; 
						        fm_size_out 	<= 14;
						        fm_depth		<= 8; // 512 todo
						        padding_out 	<= 0; 
			            	end
			            3: 
			            	begin 
			            		layer_type	<= 1; // conv
			        			activation	<= 1;

			        			fm_size		<= 14;
						        fm_depth	<= 8;  // 512 todo
						        fm_size_out <= 14; // including padding
						        padding_out <= 1;

						        kernel_num  <= 8; // 512 todo
						        kernel_size <= 3;

						        kernel_num_count <= 8 - `PARA_KERNEL*2; // 8 - `PARA_KERNEL*2 = 4 // 512 - `PARA_KERNEL*2 = 508 todo
						        write_weight_num <= (72+`PARA_Y-1)/`PARA_Y; //  3*3 * 8 = 72 // (4608+`PARA_Y-1)/`PARA_Y; 3*3 * 512 = 4608
						        next_write_weight_num <= 392; //  7*7 * 8  = 392 // 7*7* 512 = 25088 // weight_total / `PARA_Y, fc: weight_total = fm_total * PARA_Y, so fm_total * PARA_Y / PARA_Y = fm_total
			            	end
			            4:
			            	begin 
			            		layer_type		<= 2; // pool
			        			pool_type		<= 0;

						        pool_win_size	<= `POOL_SIZE;

						        fm_size 		<= 14; 
						        fm_size_out 	<= 7;
						        fm_depth		<= 8; // 512 todo
						        padding_out 	<= 0; 
			            	end
			            5:
			            	begin
			            		layer_type		<= 3; // fc
						        pre_layer_type	<= 2;

						        fm_size			<= 7;
						        fm_depth		<= 8; // 512 todo
						        fm_total_size	<= 392;// 7*7 * 8 = 392 // 7*7 * 512 = 25088

						        kernel_num		<= 16; // out put fm size, 1*1*kernel_num // 4096
						        kernel_size		<= 392; // the total size of fm
						        
						        fm_size_out 	<= 16; // 4096

						        kernel_num_count <= 16 - `PARA_Y*`PARA_KERNEL*2; // 4096 - `PARA_Y*`PARA_KERNEL*2
						        write_weight_num <= (392+`PARA_Y-1)/`PARA_Y; //  7*7 * 8 = 392 // (25088+`PARA_Y-1)/`PARA_Y; 7*7* 512 = 25088
						        next_write_weight_num <= 0; // next layer is done
			            	end
			            6:
			            	begin
			            		layer_type	<= 9; // done
			            	end
			        endcase
				end
			end
		end
	end
endmodule
