// nh means neighbourhood
`define POOL_OUT_WIDTH 16
`define NN_WIDTH 16
//`NN_WIDTH*9
`define NH_VECTOR_WIDTH 144

`define NEIGHBORHOOD_SIZE 3