module mem_controller(
);

endmodule