`define CTRL_WIDTH   30
`define SRC_2_BIAS 1