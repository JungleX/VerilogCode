// data
`define DATA_WIDTH           16       // 16 bits float