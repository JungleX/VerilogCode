// nh means neighbourhood
`define POOL_OUT_WIDTH 8
`define NN_WIDTH 8
`define NH_VECTOR_WIDTH `NN_WIDTH*9

`define NEIGHBORHOOD_SIZE 3