`define NH_VECTOR_BITWIDTH 7
`define POOL_OUT_BITWIDTH 7

`define RECT_IN_BITWIDTH 7
`define RECT_OUT_BITWIDTH 7
`define RECT_OUT_WIDTH 8

`define POOL_OUT_BITWIDTH 7
`define POOL_OUT_WIDTH 8
`define NN_BITWIDTH 7
`define NN_WIDTH 8
`define NH_VECTOR_BITWIDTH 71            //`NN_WIDTH*9-1

`define NEIGHBORHOOD_SIZE 3