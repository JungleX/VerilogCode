// nh means neighbourhood
`define POOL_OUT_WIDTH 16
`define NN_WIDTH 16
//`NN_WIDTH*9
`define NH_VECTOR_WIDTH 144

`define NEIGHBORHOOD_SIZE 3

`define POOL_WIDTH_1  55
`define POOL_HEIGHT_1 55
`define POOL_DEEP_1   96

`define POOL_WIDTH_2  27
`define POOL_HEIGHT_2 27
`define POOL_DEEP_2   256

`define POOL_WIDTH_5  13
`define POOL_HEIGHT_5 13
`define POOL_DEEP_5   256

`define COMPARE_RESULT_WIDTH 7