module dnn_accelerator(
);

mem_controller_top mem_ctrl_top();

endmodule