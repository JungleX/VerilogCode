`timescale 1ns/1ps

module top_tb();

localparam TYPE                  = "PU";
localparam integer NUM_PE        = 4;
localparam integer DATA_WIDTH    = 16;



endmodule
