`define PRECISION_OP 16
`define PRECISION_ACC 16
`define PRECISION_FRAC 8
`define num_pe 4
`define max_layers 8
