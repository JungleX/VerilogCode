0000000000000000
0000000000000001
0000000000000010
0000000000000011
0000000000000100
0000000000000101
0000000000000110
0000000000000111
0000000000001000
0000000000001001
0000000000001010
0000000000001011
0000000000001100
0000000000001101
0000000000001110
0000000000001111
0000000000010000
0000000000010001
0000000000010010
0000000000010011
0000000000010100
0000000000010101
0000000000010110
0000000000010111
0000000000011000
0000000000011001
0000000000011010
0000000000011011
0000000000011100
0000000000011101
0000000000011110
0000000000011111
0000000000100000
0000000000100001
0000000000100010
0000000000100011
0000000000100100
0000000000100101
0000000000100110
0000000000100111
0000000000101000
0000000000101001
0000000000101010
0000000000101011
0000000000101100
0000000000101101
0000000000101110
0000000000101111
0000000000110000
0000000000110001
0000000000110010
0000000000110011
0000000000110100
0000000000110101
0000000000110110
0000000000110111
0000000000111000
0000000000111001
0000000000111010
0000000000111011
0000000000111100
0000000000111101
0000000000111110
0000000000111111
0000000001000000
0000000001000001
0000000001000010
0000000001000011
0000000001000100
0000000001000101
0000000001000110
0000000001000111
0000000001001000
0000000001001001
0000000001001010
0000000001001011
0000000001001100
0000000001001101
0000000001001110
0000000001001111
0000000001010000
0000000001010001
0000000001010010
0000000001010011
0000000001010100
0000000001010101
0000000001010110
0000000001010111
0000000001011000
0000000001011001
0000000001011010
0000000001011011
0000000001011100
0000000001011101
0000000001011110
0000000001011111
0000000001100000
0000000001100001
0000000001100010
0000000001100011
0000000001100100
0000000001100101
0000000001100110
0000000001100111
0000000001101000
0000000001101001
0000000001101010
0000000001101011
0000000001101100
0000000001101101
0000000001101110
0000000001101111
0000000001110000
0000000001110001
0000000001110010
0000000001110011
0000000001110100
0000000001110101
0000000001110110
0000000001110111
0000000001111000
0000000001111001
0000000001111010
0000000001111011
0000000001111100
0000000001111101
0000000001111110
0000000001111111
0000000010000000
0000000010000001
0000000010000010
0000000010000011
0000000010000100
0000000010000101
0000000010000110
0000000010000111
0000000010001000
0000000010001001
0000000010001010
0000000010001011
0000000010001100
0000000010001101
0000000010001110
0000000010001111
0000000010010000
0000000010010001
0000000010010010
0000000010010011
0000000010010100
0000000010010101
0000000010010110
0000000010010111
0000000010011000
0000000010011001
0000000010011010
0000000010011011
0000000010011100
0000000010011101
0000000010011110
0000000010011111
0000000010100000
0000000010100001
0000000010100010
0000000010100011
0000000010100100
0000000010100101
0000000010100110
0000000010100111
0000000010101000
0000000010101001
0000000010101010
0000000010101011
0000000010101100
0000000010101101
0000000010101110
0000000010101111
0000000010110000
0000000010110001
0000000010110010
0000000010110011
0000000010110100
0000000010110101
0000000010110110
0000000010110111
0000000010111000
0000000010111001
0000000010111010
0000000010111011
0000000010111100
0000000010111101
0000000010111110
0000000010111111
0000000011000000
0000000011000001
0000000011000010
0000000011000011
0000000011000100
0000000011000101
0000000011000110
0000000011000111
0000000011001000
0000000011001001
0000000011001010
0000000011001011
0000000011001100
0000000011001101
0000000011001110
0000000011001111
0000000011010000
0000000011010001
0000000011010010
0000000011010011
0000000011010100
0000000011010101
0000000011010110
0000000011010111
0000000011011000
0000000011011001
0000000011011010
0000000011011011
0000000011011100
0000000011011101
0000000011011110
0000000011011111
0000000011100000
0000000011100001
0000000011100010
0000000011100011
0000000011100100
0000000011100101
0000000011100110
0000000011100111
0000000011101000
0000000011101001
0000000011101010
0000000011101011
0000000011101100
0000000011101101
0000000011101110
0000000011101111
0000000011110000
0000000011110001
0000000011110010
0000000011110011
0000000011110100
0000000011110101
0000000011110110
0000000011110111
0000000011111000
0000000011111001
0000000011111010
0000000011111011
0000000011111100
0000000011111101
0000000011111110
0000000011111111
0000000100000000
0000000100000001
0000000100000010
0000000100000011
0000000100000100
0000000100000101
0000000100000110
0000000100000111
0000000100001000
0000000100001001
0000000100001010
0000000100001011
0000000100001100
0000000100001101
0000000100001110
0000000100001111
0000000100010000
0000000100010001
0000000100010010
0000000100010011
0000000100010100
0000000100010101
0000000100010110
0000000100010111
0000000100011000
0000000100011001
0000000100011010
0000000100011011
0000000100011100
0000000100011101
0000000100011110
0000000100011111
0000000100100000
0000000100100001
0000000100100010
0000000100100011
0000000100100100
0000000100100101
0000000100100110
0000000100100111
0000000100101000
0000000100101001
0000000100101010
0000000100101011
0000000100101100
0000000100101101
0000000100101110
0000000100101111
0000000100110000
0000000100110001
0000000100110010
0000000100110011
0000000100110100
0000000100110101
0000000100110110
0000000100110111
0000000100111000
0000000100111001
0000000100111010
0000000100111011
0000000100111100
0000000100111101
0000000100111110
0000000100111111
0000000101000000
0000000101000001
0000000101000010
0000000101000011
0000000101000100
0000000101000101
0000000101000110
0000000101000111
0000000101001000
0000000101001001
0000000101001010
0000000101001011
0000000101001100
0000000101001101
0000000101001110
0000000101001111
0000000101010000
0000000101010001
0000000101010010
0000000101010011
0000000101010100
0000000101010101
0000000101010110
0000000101010111
0000000101011000
0000000101011001
0000000101011010
0000000101011011
0000000101011100
0000000101011101
0000000101011110
0000000101011111
0000000101100000
0000000101100001
0000000101100010
0000000101100011
0000000101100100
0000000101100101
0000000101100110
0000000101100111
0000000101101000
0000000101101001
0000000101101010
0000000101101011
0000000101101100
0000000101101101
0000000101101110
0000000101101111
0000000101110000
0000000101110001
0000000101110010
0000000101110011
0000000101110100
0000000101110101
0000000101110110
0000000101110111
0000000101111000
0000000101111001
0000000101111010
0000000101111011
0000000101111100
0000000101111101
0000000101111110
0000000101111111
0000000110000000
0000000110000001
0000000110000010
0000000110000011
0000000110000100
0000000110000101
0000000110000110
0000000110000111
0000000110001000
0000000110001001
0000000110001010
0000000110001011
0000000110001100
0000000110001101
0000000110001110
0000000110001111
0000000110010000
0000000110010001
0000000110010010
0000000110010011
0000000110010100
0000000110010101
0000000110010110
0000000110010111
0000000110011000
0000000110011001
0000000110011010
0000000110011011
0000000110011100
0000000110011101
0000000110011110
0000000110011111
0000000110100000
0000000110100001
0000000110100010
0000000110100011
0000000110100100
0000000110100101
0000000110100110
0000000110100111
0000000110101000
0000000110101001
0000000110101010
0000000110101011
0000000110101100
0000000110101101
0000000110101110
0000000110101111
0000000110110000
0000000110110001
0000000110110010
0000000110110011
0000000110110100
0000000110110101
0000000110110110
0000000110110111
0000000110111000
0000000110111001
0000000110111010
0000000110111011
0000000110111100
0000000110111101
0000000110111110
0000000110111111
0000000111000000
0000000111000001
0000000111000010
0000000111000011
0000000111000100
0000000111000101
0000000111000110
0000000111000111
0000000111001000
0000000111001001
0000000111001010
0000000111001011
0000000111001100
0000000111001101
0000000111001110
0000000111001111
0000000111010000
0000000111010001
0000000111010010
0000000111010011
0000000111010100
0000000111010101
0000000111010110
0000000111010111
0000000111011000
0000000111011001
0000000111011010
0000000111011011
0000000111011100
0000000111011101
0000000111011110
0000000111011111
0000000111100000
0000000111100001
0000000111100010
0000000111100011
0000000111100100
0000000111100101
0000000111100110
0000000111100111
0000000111101000
0000000111101001
0000000111101010
0000000111101011
0000000111101100
0000000111101101
0000000111101110
0000000111101111
0000000111110000
0000000111110001
0000000111110010
0000000111110011
0000000111110100
0000000111110101
0000000111110110
0000000111110111
0000000111111000
0000000111111001
0000000111111010
0000000111111011
0000000111111100
0000000111111101
0000000111111110
0000000111111111
0000001000000000
0000001000000001
0000001000000010
0000001000000011
0000001000000100
0000001000000101
0000001000000110
0000001000000111
0000001000001000
0000001000001001
0000001000001010
0000001000001011
0000001000001100
0000001000001101
0000001000001110
0000001000001111
0000001000010000
0000001000010001
0000001000010010
0000001000010011
0000001000010100
0000001000010101
0000001000010110
0000001000010111
0000001000011000
0000001000011001
0000001000011010
0000001000011011
0000001000011100
0000001000011101
0000001000011110
0000001000011111
0000001000100000
0000001000100001
0000001000100010
0000001000100011
0000001000100100
0000001000100101
0000001000100110
0000001000100111
0000001000101000
0000001000101001
0000001000101010
0000001000101011
0000001000101100
0000001000101101
0000001000101110
0000001000101111
0000001000110000
0000001000110001
0000001000110010
0000001000110011
0000001000110100
0000001000110101
0000001000110110
0000001000110111
0000001000111000
0000001000111001
0000001000111010
0000001000111011
0000001000111100
0000001000111101
0000001000111110
0000001000111111
0000001001000000
0000001001000001
0000001001000010
0000001001000011
0000001001000100
0000001001000101
0000001001000110
0000001001000111
0000001001001000
0000001001001001
0000001001001010
0000001001001011
0000001001001100
0000001001001101
0000001001001110
0000001001001111
0000001001010000
0000001001010001
0000001001010010
0000001001010011
0000001001010100
0000001001010101
0000001001010110
0000001001010111
0000001001011000
0000001001011001
0000001001011010
0000001001011011
0000001001011100
0000001001011101
0000001001011110
0000001001011111
0000001001100000
0000001001100001
0000001001100010
0000001001100011
0000001001100100
0000001001100101
0000001001100110
0000001001100111
0000001001101000
0000001001101001
0000001001101010
0000001001101011
0000001001101100
0000001001101101
0000001001101110
0000001001101111
0000001001110000
0000001001110001
0000001001110010
0000001001110011
0000001001110100
0000001001110101
0000001001110110
0000001001110111
0000001001111000
0000001001111001
0000001001111010
0000001001111011
0000001001111100
0000001001111101
0000001001111110
0000001001111111
0000001010000000
0000001010000001
0000001010000010
0000001010000011
0000001010000100
0000001010000101
0000001010000110
0000001010000111
0000001010001000
0000001010001001
0000001010001010
0000001010001011
0000001010001100
0000001010001101
0000001010001110
0000001010001111
0000001010010000
0000001010010001
0000001010010010
0000001010010011
0000001010010100
0000001010010101
0000001010010110
0000001010010111
0000001010011000
0000001010011001
0000001010011010
0000001010011011
0000001010011100
0000001010011101
0000001010011110
0000001010011111
0000001010100000
0000001010100001
0000001010100010
0000001010100011
0000001010100100
0000001010100101
0000001010100110
0000001010100111
0000001010101000
0000001010101001
0000001010101010
0000001010101011
0000001010101100
0000001010101101
0000001010101110
0000001010101111
0000001010110000
0000001010110001
0000001010110010
0000001010110011
0000001010110100
0000001010110101
0000001010110110
0000001010110111
0000001010111000
0000001010111001
0000001010111010
0000001010111011
0000001010111100
0000001010111101
0000001010111110
0000001010111111
0000001011000000
0000001011000001
0000001011000010
0000001011000011
0000001011000100
0000001011000101
0000001011000110
0000001011000111
0000001011001000
0000001011001001
0000001011001010
0000001011001011
0000001011001100
0000001011001101
0000001011001110
0000001011001111
0000001011010000
0000001011010001
0000001011010010
0000001011010011
0000001011010100
0000001011010101
0000001011010110
0000001011010111
0000001011011000
0000001011011001
0000001011011010
0000001011011011
0000001011011100
0000001011011101
0000001011011110
0000001011011111
0000001011100000
0000001011100001
0000001011100010
0000001011100011
0000001011100100
0000001011100101
0000001011100110
0000001011100111
0000001011101000
0000001011101001
0000001011101010
0000001011101011
0000001011101100
0000001011101101
0000001011101110
0000001011101111
0000001011110000
0000001011110001
0000001011110010
0000001011110011
0000001011110100
0000001011110101
0000001011110110
0000001011110111
0000001011111000
0000001011111001
0000001011111010
0000001011111011
0000001011111100
0000001011111101
0000001011111110
0000001011111111
0000001100000000
0000001100000001
0000001100000010
0000001100000011
0000001100000100
0000001100000101
0000001100000110
0000001100000111
0000001100001000
0000001100001001
0000001100001010
0000001100001011
0000001100001100
0000001100001101
0000001100001110
0000001100001111
0000001100010000
0000001100010001
0000001100010010
0000001100010011
0000001100010100
0000001100010101
0000001100010110
0000001100010111
0000001100011000
0000001100011001
0000001100011010
0000001100011011
0000001100011100
0000001100011101
0000001100011110
0000001100011111
0000001100100000
0000001100100001
0000001100100010
0000001100100011
0000001100100100
0000001100100101
0000001100100110
0000001100100111
0000001100101000
0000001100101001
0000001100101010
0000001100101011
0000001100101100
0000001100101101
0000001100101110
0000001100101111
0000001100110000
0000001100110001
0000001100110010
0000001100110011
0000001100110100
0000001100110101
0000001100110110
0000001100110111
0000001100111000
0000001100111001
0000001100111010
0000001100111011
0000001100111100
0000001100111101
0000001100111110
0000001100111111
0000001101000000
0000001101000001
0000001101000010
0000001101000011
0000001101000100
0000001101000101
0000001101000110
0000001101000111
0000001101001000
0000001101001001
0000001101001010
0000001101001011
0000001101001100
0000001101001101
0000001101001110
0000001101001111
0000001101010000
0000001101010001
0000001101010010
0000001101010011
0000001101010100
0000001101010101
0000001101010110
0000001101010111
0000001101011000
0000001101011001
0000001101011010
0000001101011011
0000001101011100
0000001101011101
0000001101011110
0000001101011111
0000001101100000
0000001101100001
0000001101100010
0000001101100011
0000001101100100
0000001101100101
0000001101100110
0000001101100111
0000001101101000
0000001101101001
0000001101101010
0000001101101011
0000001101101100
0000001101101101
0000001101101110
0000001101101111
0000001101110000
0000001101110001
0000001101110010
0000001101110011
0000001101110100
0000001101110101
0000001101110110
0000001101110111
0000001101111000
0000001101111001
0000001101111010
0000001101111011
0000001101111100
0000001101111101
0000001101111110
0000001101111111
0000001110000000
0000001110000001
0000001110000010
0000001110000011
0000001110000100
0000001110000101
0000001110000110
0000001110000111
0000001110001000
0000001110001001
0000001110001010
0000001110001011
0000001110001100
0000001110001101
0000001110001110
0000001110001111
0000001110010000
0000001110010001
0000001110010010
0000001110010011
0000001110010100
0000001110010101
0000001110010110
0000001110010111
0000001110011000
0000001110011001
0000001110011010
0000001110011011
0000001110011100
0000001110011101
0000001110011110
0000001110011111
0000001110100000
0000001110100001
0000001110100010
0000001110100011
0000001110100100
0000001110100101
0000001110100110
0000001110100111
0000001110101000
0000001110101001
0000001110101010
0000001110101011
0000001110101100
0000001110101101
0000001110101110
0000001110101111
0000001110110000
0000001110110001
0000001110110010
0000001110110011
0000001110110100
0000001110110101
0000001110110110
0000001110110111
0000001110111000
0000001110111001
0000001110111010
0000001110111011
0000001110111100
0000001110111101
0000001110111110
0000001110111111
0000001111000000
0000001111000001
0000001111000010
0000001111000011
0000001111000100
0000001111000101
0000001111000110
0000001111000111
0000001111001000
0000001111001001
0000001111001010
0000001111001011
0000001111001100
0000001111001101
0000001111001110
0000001111001111
0000001111010000
0000001111010001
0000001111010010
0000001111010011
0000001111010100
0000001111010101
0000001111010110
0000001111010111
0000001111011000
0000001111011001
0000001111011010
0000001111011011
0000001111011100
0000001111011101
0000001111011110
0000001111011111
0000001111100000
0000001111100001
0000001111100010
0000001111100011
0000001111100100
0000001111100101
0000001111100110
0000001111100111
0000001111101000
0000001111101001
0000001111101010
0000001111101011
0000001111101100
0000001111101101
0000001111101110
0000001111101111
0000001111110000
0000001111110001
0000001111110010
0000001111110011
0000001111110100
0000001111110101
0000001111110110
0000001111110111
0000001111111000
0000001111111001
0000001111111010
0000001111111011
0000001111111100
0000001111111101
0000001111111110
0000001111111111
0000010000000000
0000010000000001
0000010000000010
0000010000000011
0000010000000100
0000010000000101
0000010000000110
0000010000000111
0000010000001000
0000010000001001
0000010000001010
0000010000001011
0000010000001100
0000010000001101
0000010000001110
0000010000001111
0000010000010000
0000010000010001
0000010000010010
0000010000010011
0000010000010100
0000010000010101
0000010000010110
0000010000010111
0000010000011000
0000010000011001
0000010000011010
0000010000011011
0000010000011100
0000010000011101
0000010000011110
0000010000011111
0000010000100000
0000010000100001
0000010000100010
0000010000100011
0000010000100100
0000010000100101
0000010000100110
0000010000100111
0000010000101000
0000010000101001
0000010000101010
0000010000101011
0000010000101100
0000010000101101
0000010000101110
0000010000101111
0000010000110000
0000010000110001
0000010000110010
0000010000110011
0000010000110100
0000010000110101
0000010000110110
0000010000110111
0000010000111000
0000010000111001
0000010000111010
0000010000111011
0000010000111100
0000010000111101
0000010000111110
0000010000111111
0000010001000000
0000010001000001
0000010001000010
0000010001000011
0000010001000100
0000010001000101
0000010001000110
0000010001000111
0000010001001000
0000010001001001
0000010001001010
0000010001001011
0000010001001100
0000010001001101
0000010001001110
0000010001001111
0000010001010000
0000010001010001
0000010001010010
0000010001010011
0000010001010100
0000010001010101
0000010001010110
0000010001010111
0000010001011000
0000010001011001
0000010001011010
0000010001011011
0000010001011100
0000010001011101
0000010001011110
0000010001011111
0000010001100000
0000010001100001
0000010001100010
0000010001100011
0000010001100100
0000010001100101
0000010001100110
0000010001100111
0000010001101000
0000010001101001
0000010001101010
0000010001101011
0000010001101100
0000010001101101
0000010001101110
0000010001101111
0000010001110000
0000010001110001
0000010001110010
0000010001110011
0000010001110100
0000010001110101
0000010001110110
0000010001110111
0000010001111000
0000010001111001
0000010001111010
0000010001111011
0000010001111100
0000010001111101
0000010001111110
0000010001111111
0000010010000000
0000010010000001
0000010010000010
0000010010000011
0000010010000100
0000010010000101
0000010010000110
0000010010000111
0000010010001000
0000010010001001
0000010010001010
0000010010001011
0000010010001100
0000010010001101
0000010010001110
0000010010001111
0000010010010000
0000010010010001
0000010010010010
0000010010010011
0000010010010100
0000010010010101
0000010010010110
0000010010010111
0000010010011000
0000010010011001
0000010010011010
0000010010011011
0000010010011100
0000010010011101
0000010010011110
0000010010011111
0000010010100000
0000010010100001
0000010010100010
0000010010100011
0000010010100100
0000010010100101
0000010010100110
0000010010100111
0000010010101000
0000010010101001
0000010010101010
0000010010101011
0000010010101100
0000010010101101
0000010010101110
0000010010101111
0000010010110000
0000010010110001
0000010010110010
0000010010110011
0000010010110100
0000010010110101
0000010010110110
0000010010110111
0000010010111000
0000010010111001
0000010010111010
0000010010111011
0000010010111100
0000010010111101
0000010010111110
0000010010111111
0000010011000000
0000010011000001
0000010011000010
0000010011000011
0000010011000100
0000010011000101
0000010011000110
0000010011000111
0000010011001000
0000010011001001
0000010011001010
0000010011001011
0000010011001100
0000010011001101
0000010011001110
0000010011001111
0000010011010000
0000010011010001
0000010011010010
0000010011010011
0000010011010100
0000010011010101
0000010011010110
0000010011010111
0000010011011000
0000010011011001
0000010011011010
0000010011011011
0000010011011100
0000010011011101
0000010011011110
0000010011011111
0000010011100000
0000010011100001
0000010011100010
0000010011100011
0000010011100100
0000010011100101
0000010011100110
0000010011100111
0000010011101000
0000010011101001
0000010011101010
0000010011101011
0000010011101100
0000010011101101
0000010011101110
0000010011101111
0000010011110000
0000010011110001
0000010011110010
0000010011110011
0000010011110100
0000010011110101
0000010011110110
0000010011110111
0000010011111000
0000010011111001
0000010011111010
0000010011111011
0000010011111100
0000010011111101
0000010011111110
0000010011111111
0000010100000000
0000010100000001
0000010100000010
0000010100000011
0000010100000100
0000010100000101
0000010100000110
0000010100000111
0000010100001000
0000010100001001
0000010100001010
0000010100001011
0000010100001100
0000010100001101
0000010100001110
0000010100001111
0000010100010000
0000010100010001
0000010100010010
0000010100010011
0000010100010100
0000010100010101
0000010100010110
0000010100010111
0000010100011000
0000010100011001
0000010100011010
0000010100011011
0000010100011100
0000010100011101
0000010100011110
0000010100011111
0000010100100000
0000010100100001
0000010100100010
0000010100100011
0000010100100100
0000010100100101
0000010100100110
0000010100100111
0000010100101000
0000010100101001
0000010100101010
0000010100101011
0000010100101100
0000010100101101
0000010100101110
0000010100101111
0000010100110000
0000010100110001
0000010100110010
0000010100110011
0000010100110100
0000010100110101
0000010100110110
0000010100110111
0000010100111000
0000010100111001
0000010100111010
0000010100111011
0000010100111100
0000010100111101
0000010100111110
0000010100111111
0000010101000000
0000010101000001
0000010101000010
0000010101000011
0000010101000100
0000010101000101
0000010101000110
0000010101000111
0000010101001000
0000010101001001
0000010101001010
0000010101001011
0000010101001100
0000010101001101
0000010101001110
0000010101001111
0000010101010000
0000010101010001
0000010101010010
0000010101010011
0000010101010100
0000010101010101
0000010101010110
0000010101010111
0000010101011000
0000010101011001
0000010101011010
0000010101011011
0000010101011100
0000010101011101
0000010101011110
0000010101011111
0000010101100000
0000010101100001
0000010101100010
0000010101100011
0000010101100100
0000010101100101
0000010101100110
0000010101100111
0000010101101000
0000010101101001
0000010101101010
0000010101101011
0000010101101100
0000010101101101
0000010101101110
0000010101101111
0000010101110000
0000010101110001
0000010101110010
0000010101110011
0000010101110100
0000010101110101
0000010101110110
0000010101110111
0000010101111000
0000010101111001
0000010101111010
0000010101111011
0000010101111100
0000010101111101
0000010101111110
0000010101111111
0000010110000000
0000010110000001
0000010110000010
0000010110000011
0000010110000100
0000010110000101
0000010110000110
0000010110000111
0000010110001000
0000010110001001
0000010110001010
0000010110001011
0000010110001100
0000010110001101
0000010110001110
0000010110001111
0000010110010000
0000010110010001
0000010110010010
0000010110010011
0000010110010100
0000010110010101
0000010110010110
0000010110010111
0000010110011000
0000010110011001
0000010110011010
0000010110011011
0000010110011100
0000010110011101
0000010110011110
0000010110011111
0000010110100000
0000010110100001
0000010110100010
0000010110100011
0000010110100100
0000010110100101
0000010110100110
0000010110100111
0000010110101000
0000010110101001
0000010110101010
0000010110101011
0000010110101100
0000010110101101
0000010110101110
0000010110101111
0000010110110000
0000010110110001
0000010110110010
0000010110110011
0000010110110100
0000010110110101
0000010110110110
0000010110110111
0000010110111000
0000010110111001
0000010110111010
0000010110111011
0000010110111100
0000010110111101
0000010110111110
0000010110111111
0000010111000000
0000010111000001
0000010111000010
0000010111000011
0000010111000100
0000010111000101
0000010111000110
0000010111000111
0000010111001000
0000010111001001
0000010111001010
0000010111001011
0000010111001100
0000010111001101
0000010111001110
0000010111001111
0000010111010000
0000010111010001
0000010111010010
0000010111010011
0000010111010100
0000010111010101
0000010111010110
0000010111010111
0000010111011000
0000010111011001
0000010111011010
0000010111011011
0000010111011100
0000010111011101
0000010111011110
0000010111011111
0000010111100000
0000010111100001
0000010111100010
0000010111100011
0000010111100100
0000010111100101
0000010111100110
0000010111100111
0000010111101000
0000010111101001
0000010111101010
0000010111101011
0000010111101100
0000010111101101
0000010111101110
0000010111101111
0000010111110000
0000010111110001
0000010111110010
0000010111110011
0000010111110100
0000010111110101
0000010111110110
0000010111110111
0000010111111000
0000010111111001
0000010111111010
0000010111111011
0000010111111100
0000010111111101
0000010111111110
0000010111111111
0000011000000000
0000011000000001
0000011000000010
0000011000000011
0000011000000100
0000011000000101
0000011000000110
0000011000000111
0000011000001000
0000011000001001
0000011000001010
0000011000001011
0000011000001100
0000011000001101
0000011000001110
0000011000001111
0000011000010000
0000011000010001
0000011000010010
0000011000010011
0000011000010100
0000011000010101
0000011000010110
0000011000010111
0000011000011000
0000011000011001
0000011000011010
0000011000011011
0000011000011100
0000011000011101
0000011000011110
0000011000011111
0000011000100000
0000011000100001
0000011000100010
0000011000100011
0000011000100100
0000011000100101
0000011000100110
0000011000100111
0000011000101000
0000011000101001
0000011000101010
0000011000101011
0000011000101100
0000011000101101
0000011000101110
0000011000101111
0000011000110000
0000011000110001
0000011000110010
0000011000110011
0000011000110100
0000011000110101
0000011000110110
0000011000110111
0000011000111000
0000011000111001
0000011000111010
0000011000111011
0000011000111100
0000011000111101
0000011000111110
0000011000111111
0000011001000000
0000011001000001
0000011001000010
0000011001000011
0000011001000100
0000011001000101
0000011001000110
0000011001000111
0000011001001000
0000011001001001
0000011001001010
0000011001001011
0000011001001100
0000011001001101
0000011001001110
0000011001001111
0000011001010000
0000011001010001
0000011001010010
0000011001010011
0000011001010100
0000011001010101
0000011001010110
0000011001010111
0000011001011000
0000011001011001
0000011001011010
0000011001011011
0000011001011100
0000011001011101
0000011001011110
0000011001011111
0000011001100000
0000011001100001
0000011001100010
0000011001100011
0000011001100100
0000011001100101
0000011001100110
0000011001100111
0000011001101000
0000011001101001
0000011001101010
0000011001101011
0000011001101100
0000011001101101
0000011001101110
0000011001101111
0000011001110000
0000011001110001
0000011001110010
0000011001110011
0000011001110100
0000011001110101
0000011001110110
0000011001110111
0000011001111000
0000011001111001
0000011001111010
0000011001111011
0000011001111100
0000011001111101
0000011001111110
0000011001111111
0000011010000000
0000011010000001
0000011010000010
0000011010000011
0000011010000100
0000011010000101
0000011010000110
0000011010000111
0000011010001000
0000011010001001
0000011010001010
0000011010001011
0000011010001100
0000011010001101
0000011010001110
0000011010001111
0000011010010000
0000011010010001
0000011010010010
0000011010010011
0000011010010100
0000011010010101
0000011010010110
0000011010010111
0000011010011000
0000011010011001
0000011010011010
0000011010011011
0000011010011100
0000011010011101
0000011010011110
0000011010011111
0000011010100000
0000011010100001
0000011010100010
0000011010100011
0000011010100100
0000011010100101
0000011010100110
0000011010100111
0000011010101000
0000011010101001
0000011010101010
0000011010101011
0000011010101100
0000011010101101
0000011010101110
0000011010101111
0000011010110000
0000011010110001
0000011010110010
0000011010110011
0000011010110100
0000011010110101
0000011010110110
0000011010110111
0000011010111000
0000011010111001
0000011010111010
0000011010111011
0000011010111100
0000011010111101
0000011010111110
0000011010111111
0000011011000000
0000011011000001
0000011011000010
0000011011000011
0000011011000100
0000011011000101
0000011011000110
0000011011000111
0000011011001000
0000011011001001
0000011011001010
0000011011001011
0000011011001100
0000011011001101
0000011011001110
0000011011001111
0000011011010000
0000011011010001
0000011011010010
0000011011010011
0000011011010100
0000011011010101
0000011011010110
0000011011010111
0000011011011000
0000011011011001
0000011011011010
0000011011011011
0000011011011100
0000011011011101
0000011011011110
0000011011011111
0000011011100000
0000011011100001
0000011011100010
0000011011100011
0000011011100100
0000011011100101
0000011011100110
0000011011100111
0000011011101000
0000011011101001
0000011011101010
0000011011101011
0000011011101100
0000011011101101
0000011011101110
0000011011101111
0000011011110000
0000011011110001
0000011011110010
0000011011110011
0000011011110100
0000011011110101
0000011011110110
0000011011110111
0000011011111000
0000011011111001
0000011011111010
0000011011111011
0000011011111100
0000011011111101
0000011011111110
0000011011111111
0000011100000000
0000011100000001
0000011100000010
0000011100000011
0000011100000100
0000011100000101
0000011100000110
0000011100000111
0000011100001000
0000011100001001
0000011100001010
0000011100001011
0000011100001100
0000011100001101
0000011100001110
0000011100001111
0000011100010000
0000011100010001
0000011100010010
0000011100010011
0000011100010100
0000011100010101
0000011100010110
0000011100010111
0000011100011000
0000011100011001
0000011100011010
0000011100011011
0000011100011100
0000011100011101
0000011100011110
0000011100011111
0000011100100000
0000011100100001
0000011100100010
0000011100100011
0000011100100100
0000011100100101
0000011100100110
0000011100100111
0000011100101000
0000011100101001
0000011100101010
0000011100101011
0000011100101100
0000011100101101
0000011100101110
0000011100101111
0000011100110000
0000011100110001
0000011100110010
0000011100110011
0000011100110100
0000011100110101
0000011100110110
0000011100110111
0000011100111000
0000011100111001
0000011100111010
0000011100111011
0000011100111100
0000011100111101
0000011100111110
0000011100111111
0000011101000000
0000011101000001
0000011101000010
0000011101000011
0000011101000100
0000011101000101
0000011101000110
0000011101000111
0000011101001000
0000011101001001
0000011101001010
0000011101001011
0000011101001100
0000011101001101
0000011101001110
0000011101001111
0000011101010000
0000011101010001
0000011101010010
0000011101010011
0000011101010100
0000011101010101
0000011101010110
0000011101010111
0000011101011000
0000011101011001
0000011101011010
0000011101011011
0000011101011100
0000011101011101
0000011101011110
0000011101011111
0000011101100000
0000011101100001
0000011101100010
0000011101100011
0000011101100100
0000011101100101
0000011101100110
0000011101100111
0000011101101000
0000011101101001
0000011101101010
0000011101101011
0000011101101100
0000011101101101
0000011101101110
0000011101101111
0000011101110000
0000011101110001
0000011101110010
0000011101110011
0000011101110100
0000011101110101
0000011101110110
0000011101110111
0000011101111000
0000011101111001
0000011101111010
0000011101111011
0000011101111100
0000011101111101
0000011101111110
0000011101111111
0000011110000000
0000011110000001
0000011110000010
0000011110000011
0000011110000100
0000011110000101
0000011110000110
0000011110000111
0000011110001000
0000011110001001
0000011110001010
0000011110001011
0000011110001100
0000011110001101
0000011110001110
0000011110001111
0000011110010000
0000011110010001
0000011110010010
0000011110010011
0000011110010100
0000011110010101
0000011110010110
0000011110010111
0000011110011000
0000011110011001
0000011110011010
0000011110011011
0000011110011100
0000011110011101
0000011110011110
0000011110011111
0000011110100000
0000011110100001
0000011110100010
0000011110100011
0000011110100100
0000011110100101
0000011110100110
0000011110100111
0000011110101000
0000011110101001
0000011110101010
0000011110101011
0000011110101100
0000011110101101
0000011110101110
0000011110101111
0000011110110000
0000011110110001
0000011110110010
0000011110110011
0000011110110100
0000011110110101
0000011110110110
0000011110110111
0000011110111000
0000011110111001
0000011110111010
0000011110111011
0000011110111100
0000011110111101
0000011110111110
0000011110111111
0000011111000000
0000011111000001
0000011111000010
0000011111000011
0000011111000100
0000011111000101
0000011111000110
0000011111000111
0000011111001000
0000011111001001
0000011111001010
0000011111001011
0000011111001100
0000011111001101
0000011111001110
0000011111001111
0000011111010000
0000011111010001
0000011111010010
0000011111010011
0000011111010100
0000011111010101
0000011111010110
0000011111010111
0000011111011000
0000011111011001
0000011111011010
0000011111011011
0000011111011100
0000011111011101
0000011111011110
0000011111011111
0000011111100000
0000011111100001
0000011111100010
0000011111100011
0000011111100100
0000011111100101
0000011111100110
0000011111100111
0000011111101000
0000011111101001
0000011111101010
0000011111101011
0000011111101100
0000011111101101
0000011111101110
0000011111101111
0000011111110000
0000011111110001
0000011111110010
0000011111110011
0000011111110100
0000011111110101
0000011111110110
0000011111110111
0000011111111000
0000011111111001
0000011111111010
0000011111111011
0000011111111100
0000011111111101
0000011111111110
0000011111111111