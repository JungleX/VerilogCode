`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: SJTU Tcloud FPGA Group
// Engineer: 
// 
// Create Date: 2017/05/26 16:53:16
// Design Name: 
// Module Name: multX11_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
//  
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`define clk_period 10

`include "alexnet_parameters.vh"

module multX11_tb();
	reg clk;
	reg rst;
    reg ena;

    reg [`CONV_MAX_LINE_SIZE - 1:0] data;     
    
    reg [`CONV_MAX_LINE_SIZE - 1:0] weight;   

    wire [`DATA_WIDTH - 1:0] out;

    multX11 conv(
    	.clk(clk),
    	.rst(rst),
    	.ena(ena),

    	.data(data),
    	.weight(weight),

    	.out(out)
    	);

    initial 
        clk = 1'b0;
    always #(`clk_period/2)clk = ~clk;


    initial begin
    	#0
    	rst = 0;

    	#(`clk_period/2)
    	ena = 1;
    	rst = 1;
    	data   = {16'b0011110000000000, 16'b0100000000000000, 16'b0100001000000000, 16'b0011110000000000, 16'b0100000000000000, 
    			  16'b0100001000000000, 16'b0011110000000000, 16'b0100000000000000, 16'b0100001000000000, 16'b0100001000000000,
    			  16'b0100000000000000};
    			 // 1,2,3,1,2,3,1,2,3,3,2
    	weight = {16'b0011110000000000, 16'b1011110000000000, 16'b0011110000000000, 16'b1011110000000000, 16'b0011110000000000, 
    	          16'b1011110000000000, 16'b0011110000000000, 16'b1011110000000000, 16'b0011110000000000, 16'b1011110000000000,
    	          16'b0011110000000000
    	      	 };
    	      	 // 1,-1,1,-1,1,-1,1,-1,1,-1,1
    	// result = 1 = 3c00;

    	#(`clk_period+`clk_period/2)
    	data   = {16'b0011110000000000, 16'b0100000000000000, 16'b0100001000000000, 16'b0011110000000000, 16'b0100000000000000, 
    			  16'b0100001000000000, 16'b0011110000000000, 16'b0100000000000000, 16'b0100001000000000, 16'b0100001000000000,
    			  16'b0011110000000000};
    			 // 1,2,3,1,2,3,1,2,3,3,1
    	weight = {16'b1011110000000000, 16'b1011110000000000, 16'b1011110000000000, 16'b1011110000000000, 16'b1011110000000000, 
    	          16'b1011110000000000, 16'b1011110000000000, 16'b1011110000000000, 16'b1011110000000000, 16'b1011110000000000,
    	          16'b1011110000000000
    	      	 };
    	      	 // -1,-1,-1,-1,-1,-1,-1,-1,-1,-1,-1
    	// result = -22 = cd80;

    	#`clk_period
    	data   = {16'b1011110000000000, 16'b1100000000000000, 16'b1100001000000000, 16'b1011110000000000, 16'b1100000000000000, 
    			  16'b1100001000000000, 16'b1011110000000000, 16'b1100000000000000, 16'b1100001000000000, 16'b1100001000000000,
    			  16'b1100000000000000};
    			 // -1,-2,-3,-1,-2,-3,-1,-2,-3,-3,-2
    	weight = {16'b0011110000000000, 16'b1011110000000000, 16'b0011110000000000, 16'b1011110000000000, 16'b0011110000000000, 
    	          16'b1011110000000000, 16'b0011110000000000, 16'b1011110000000000, 16'b0011110000000000, 16'b1011110000000000,
    	          16'b0011110000000000
    	      	 };
    	      	 // 1,-1,1,-1,1,-1,1,-1,1,-1,1
    	// result = -1 = bc00;

    	#`clk_period
    	data   = 0;
    	weight = 0;

    	#(`clk_period*9)
    	rst = 0;

    end

endmodule
