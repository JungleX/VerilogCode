`define SRC_2_BIAS 1