`include "common.vh"

module PE
(
    input wire              clk,
    input wire              reset,
    input wire [ `CTRL_WIDTH - 1 : 0 ]              ctrl
);

endmodule