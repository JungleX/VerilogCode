module mem_controller_top(
);

mem_controller u_mem_ctrl(
);

endmodule